** Profile: "SCHEMATIC1-bias"  [ c:\users\taylorrc\documents\testingcircuit-pspicefiles\schematic1\bias.sim ] 

** Creating circuit file "bias.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Cadence/SPB_16.6/tools/pspice/library/irf.lib" 
.LIB "C:/Cadence/SPB_16.6/tools/pspice/library/opamp.lib" 
.LIB "C:/Cadence/SPB_16.6/tools/pspice/library/ebipolar.lib" 
.LIB "C:/Cadence/RHIT_Libraries/RHIT_Libraries/Class.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 180 0 0.01 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
